package GeneralVariables;

parameter DATA_WIDTH = 31;

endpackage