package GeneralVariables;

  parameter logic[5:0] DATA_WIDTH = 31;

endpackage
